���      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.1.3�ub�n_estimators�K�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h)�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Age��Sex��ChestPainType��	RestingBP��Cholesterol��	FastingBS��
RestingECG�et�b�n_features_in_�K�
n_outputs_�K�classes_�h(h+K ��h-��R�(KK��h2�i4�����R�(K�<�NNNJ����J����K t�b�C       �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh$hNhJ�
hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h2�f8�����R�(KhKNNNJ����J����K t�b�C              �?�t�bhOh&�scalar���h2�i8�����R�(KhKNNNJ����J����K t�bC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hK�
node_count�Ky�nodes�h(h+K ��h-��R�(KKy��h2�V56�����R�(Kh6N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hhcK ��h�hcK��h�hcK��h�h[K��h�h[K ��h�hcK(��h�h[K0��uK8KKt�b�Bx         f                    @K@�`��ie�?�           ��@                          Ph@������?�            `w@                           �C@|�n��T�?F            @[@                           �?���N8�?             5@                          �`@r�q��?             2@       	                    @A@���!pc�?	             &@                           �?      �?              @������������������������       �                     �?������������������������       �                     �?
                           �?�<ݚ�?             "@������������������������       �                      @������������������������       �                     @������������������������       �                     @                            B@�q�q�?             @������������������������       �                     �?������������������������       �                      @                          Pf@����!p�?7             V@                           �?����p�?+             Q@������������������������       �                     @������������������������       �        '            �O@������������������������       �                     4@       [                    �?���	��?�            �p@       (                    @F@�9+�Q�?�             m@                           �?�p ��?3            �T@                           �?     ��?             @@������������������������       �                     @������������������������       �                     =@                          �h@j�q����?!             I@������������������������       �                     @       !                   �k@��E�B��?             �G@                            �?     ��?	             0@������������������������       �                     @������������������������       �                     &@"       '                    �?�g�y��?             ?@#       $                    @D@�X�<ݺ?             2@������������������������       �                      @%       &                   �_@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     *@)       B                    �?�w��#��?b            �b@*       ?                    �?<�A+K&�?/             S@+       6                    �?r�q��?+             R@,       5                   p@؇���X�?             5@-       .                    �F@�q�q�?             "@������������������������       �                      @/       0                   m@և���X�?             @������������������������       �                     @1       4                   o@      �?             @2       3                     H@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@7       <                   �p@@�0�!��?             �I@8       ;                    @H@P���Q�?             D@9       :                    �?�<ݚ�?             "@������������������������       �                      @������������������������       �                     @������������������������       �                     ?@=       >                    �?���|���?             &@������������������������       �                     @������������������������       �                     @@       A                    �?      �?             @������������������������       �                     �?������������������������       �                     @C       P                   �p@��+��?3            �R@D       M                    @J@
j*D>�?#             J@E       H                   �o@      �?             E@F       G                    �?����e��?            �@@������������������������       �                     4@������������������������       �        
             *@I       L                   @p@�����H�?             "@J       K                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @N       O                    �?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@Q       V                   Hs@���!pc�?             6@R       U                    �?     ��?             0@S       T                    �?      �?	             (@������������������������       �                     "@������������������������       �                     @������������������������       �                     @W       X                    @J@      �?             @������������������������       �                     �?Y       Z                    �?���Q��?             @������������������������       �                     @������������������������       �                      @\       c                    �J@�eP*L��?            �@@]       `                    �?��}*_��?             ;@^       _                    �?�r����?             .@������������������������       �                      @������������������������       �        
             *@a       b                    �?�q�q�?             (@������������������������       �                      @������������������������       �                     @d       e                   �b@r�q��?             @������������������������       �                     @������������������������       �                     �?g       r                   u@DG��L�?�            �v@h       k                   Xr@'Ko���?�            @u@i       j                    �?�luL3�?�            Ps@������������������������       �                     ?@������������������������       �        �            `q@l       o                   Ps@f���M�?             ?@m       n                    �?      �?             2@������������������������       �                     "@������������������������       �                     "@p       q                     L@8�Z$���?             *@������������������������       �                      @������������������������       �                     &@s       t                   ``@z�G�z�?             4@������������������������       �                      @u       v                   �`@�q�q�?             (@������������������������       �                     @w       x                   Hx@�����H�?             "@������������������������       �                     �?������������������������       �                      @�t�b�values�h(h+K ��h-��R�(KKyKK��h[�B�       @b@     `�@      V@     �q@      $@     �X@      @      0@      @      .@      @       @      �?      �?      �?                      �?       @      @       @                      @              @       @      �?              �?       @              @     �T@      @     �O@      @                     �O@              4@     �S@     `g@     �O@      e@      (@     �Q@      @      =@      @                      =@      "@     �D@      @              @     �D@      @      &@      @                      &@      �?      >@      �?      1@               @      �?      "@              "@      �?                      *@     �I@     �X@      *@     �O@      (@      N@      @      2@      @      @               @      @      @              @      @      �?       @      �?       @                      �?      �?                      (@      "@      E@       @      C@       @      @       @                      @              ?@      @      @      @                      @      �?      @      �?                      @      C@      B@      6@      >@      5@      5@      4@      *@      4@                      *@      �?       @      �?      @      �?                      @              @      �?      "@      �?                      "@      0@      @      *@      @      "@      @      "@                      @      @              @      @              �?      @       @      @                       @      .@      2@      $@      1@       @      *@       @                      *@       @      @       @                      @      @      �?      @                      �?      M@     �r@      E@     �r@      ?@     `q@      ?@                     `q@      &@      4@      "@      "@      "@                      "@       @      &@       @                      &@      0@      @       @               @      @              @       @      �?              �?       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ/��hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvK/hwh(h+K ��h-��R�(KK/��h~�BH
         $                    �?>�y@��?�           ��@                           �@@(�.���?�            0x@                            @@�q�q�?             @������������������������       �                     �?������������������������       �                      @       !                    �?     ��?�             x@                           �?���|��?�            �r@                          pw@�>4և��?�             l@	       
                    �?�uX��?�             k@������������������������       �                    �@@������������������������       �        r             g@������������������������       �                     @                           �l@��(�2Y�?+            �R@                          `k@�S����?             �L@                          @W@0��_��?            �J@                          `X@X�EQ]N�?            �E@                           @N@����X�?             @������������������������       �                     @������������������������       �                      @                          �b@�8��8��?             B@                           �I@�FVQ&�?            �@@                           �?8�Z$���?             *@������������������������       �                      @������������������������       �                     &@������������������������       �                     4@                          Pd@�q�q�?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@������������������������       �                     @������������������������       �                     1@"       #                    �?���1j	�?<            �U@������������������������       �                     @������������������������       �        7            @T@%       ,                   �Z@�`�����?�            �u@&       '                   �c@p�ݯ��?             3@������������������������       �                     @(       )                    @H@؇���X�?             ,@������������������������       �                     "@*       +                    �?���Q��?             @������������������������       �                     @������������������������       �                      @-       .                    �?�yQ�|�?�            �t@������������������������       �        9            �V@������������������������       �        �            �m@�t�bh�h(h+K ��h-��R�(KK/KK��h[�B�       �c@      �@      L@     �t@       @      �?              �?       @              K@     �t@     �H@      o@      D@      g@     �@@      g@     �@@                      g@      @              "@     @P@      "@      H@      @      H@      @      C@       @      @              @       @              @     �@@       @      ?@       @      &@       @                      &@              4@      �?       @      �?      �?      �?                      �?              �?              $@      @                      1@      @     @T@      @                     @T@     �Y@     �n@      (@      @              @      (@       @      "@              @       @      @                       @     �V@     �m@     �V@                     �m@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJu�7hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvKhwh(h+K ��h-��R�(KK��h~�B                            �^@ ���wJ�?�           ��@                          �[@j[j�v��?�            �l@                           �?L� P?)�??            @X@������������������������       �                     3@������������������������       �        2            �S@       	                     D@�X���?Y            �`@                           �?�8��8��?             8@������������������������       �                      @������������������������       �                     6@
                           �?���B��?I             [@������������������������       �                    �E@������������������������       �        4            @P@                          �_@䩱��<�?G           �@                           �?P�Lt�<�?             C@������������������������       �                     @@                           �?r�q��?             @������������������������       �                     @                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �?@	*�+�?,           0}@������������������������       �        4             T@������������������������       �        �            0x@�t�bh�h(h+K ��h-��R�(KKKK��h[�Bp        b@     h�@      P@     �d@      3@     �S@      3@                     �S@     �F@     �U@       @      6@       @                      6@     �E@     @P@     �E@                     @P@     @T@     �z@      �?     �B@              @@      �?      @              @      �?       @      �?                       @      T@     0x@      T@                     0x@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��!XhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvK#hwh(h+K ��h-��R�(KK#��h~�B�                             �a@�Z{����?�           ��@                          @^@�:�]��?c             c@                           �?*
;&���?             G@������������������������       �                     1@                           �?>���Rp�?             =@                            K@���B���?             :@                           @B@�q�q�?             (@������������������������       �                     @	       
                    �?X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @                          `X@@4և���?	             ,@                           @N@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     &@                            K@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           I@�f�¦ζ?D            �Z@                           �Q@�X�<ݺ?:            �V@                           @I@`��F:u�?8            �U@                           �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @                           �?�g<a�?2            @S@������������������������       �                      @������������������������       �        0            �R@                           `R@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        
             1@!       "                    �?T��L�?|           (�@������������������������       �        a            �b@������������������������       �                   {@�t�bh�h(h+K ��h-��R�(KK#KK��h[�B0        d@     ��@      (@     �a@      @     �C@              1@      @      6@      @      5@      @       @              @      @      @      @                      @      �?      *@      �?       @               @      �?                      &@       @      �?              �?       @              @     �Y@      @     @U@      @     �T@       @       @       @                       @       @     �R@       @                     �R@      �?       @      �?                       @              1@     �b@     {@     �b@                     {@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJC�NhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvK-hwh(h+K ��h-��R�(KK-��h~�B�	         
                    �?6_1����?�           ��@                          pv@�MG��?           ��@                           �?:=G���?t            �@������������������������       �        P            �_@������������������������       �        $           `z@                           �?ҳ�wY;�?             1@������������������������       �                     "@       	                    b@      �?              @������������������������       �                     @������������������������       �                      @                           @@@Р�31�?d             e@������������������������       �                     @                          �i@p���I�?c            �d@                           �?`<)�+�?-            @S@                           S@P����?"            �M@                           �?�Ń��̧?             E@������������������������       �        
             3@                           _@�nkK�?             7@                           �?      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     .@������������������������       �        	             1@                           @�����H�?             2@                            Q@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?                          @_@r�q��?             @������������������������       �                     �?������������������������       �                     @       $                    @L@��f��?6            @V@        !                   �i@�	j*D�?             J@������������������������       �                     @"       #                    �?      �?             H@������������������������       �                     (@������������������������       �                     B@%       ,                   �`@@-�_ .�?            �B@&       +                    �?r�q��?             (@'       (                   (p@�C��2(�?             &@������������������������       �                      @)       *                     O@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     9@�t�bh�h(h+K ��h-��R�(KK-KK��h[�B�        d@     �@      a@     �z@     �_@     `z@     �_@                     `z@      &@      @      "@               @      @              @       @              8@      b@      @              5@      b@      @     �R@      �?      M@      �?     �D@              3@      �?      6@      �?      @      �?                      @              .@              1@       @      0@      �?      &@              &@      �?              �?      @      �?                      @      2@     �Q@      0@      B@      @              (@      B@      (@                      B@       @     �A@       @      $@      �?      $@               @      �?       @      �?                       @      �?                      9@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�R�[hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvKhwh(h+K ��h-��R�(KK��h~�C�                           �?>�y@��?�           ��@������������������������       �        f            �c@������������������������       �        g            �@�t�bh�h(h+K ��h-��R�(KKKK��h[�C0     �c@      �@     �c@                      �@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�v}hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvKhwh(h+K ��h-��R�(KK��h~�C�                           �?H�ig��?�           ��@������������������������       �        g             e@������������������������       �        f           ��@�t�bh�h(h+K ��h-��R�(KKKK��h[�C0      e@     ��@      e@                     ��@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJg}�XhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKǅ�h~�B�+         �                    �?�M�dt��?�           ��@       �                   Xr@0�����?{           H�@       8                    �?L�zF�?K           �@       7                   Hq@ףp=
�?�            @p@       2                    �N@�Ӆ�0�?�            `m@       '                    @K@T�\�9�?w             g@       $                   �p@�̐d��?G            @Z@       #                   `a@���2j��?E            �Y@	                           �?2%ޑ��?/            �Q@
                          �`@������?	             .@                           �?8�Z$���?             *@������������������������       �                      @������������������������       �                     &@������������������������       �                      @                          @[@X�;�^o�?&            �K@                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �?4��?�?$             J@                           j@@4և���?             E@                          pi@      �?             8@                           �?���}<S�?             7@������������������������       �                      @������������������������       �                     5@������������������������       �                     �?������������������������       �                     2@                            �G@z�G�z�?             $@                           @F@      �?              @                          �j@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @!       "                   �^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @@%       &                   ``@�q�q�?             @������������������������       �                     �?������������������������       �                      @(       )                   `i@x�G�z�?0             T@������������������������       �                     <@*       +                   �i@0G���ջ?             J@������������������������       �                     �?,       -                    �?`'�J�?            �I@������������������������       �                     ,@.       /                    @L@@-�_ .�?            �B@������������������������       �                     2@0       1                    �?�KM�]�?             3@������������������������       �                      @������������������������       �                     1@3       6                   �p@z�G�z�?             I@4       5                    �?��0{9�?            �G@������������������������       �                     @������������������������       �                     D@������������������������       �                     @������������������������       �                     9@9       R                   h@@�j���?�            @o@:       G                    @O@0��_��?'            �J@;       F                    �? �#�Ѵ�?            �E@<       =                   a@�}�+r��?             C@������������������������       �        	             &@>       E                    �F@�>����?             ;@?       @                    �C@z�G�z�?             $@������������������������       �                     @A       B                   �\@      �?             @������������������������       �                     �?C       D                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        
             1@������������������������       �                     @H       I                    �?�z�G��?             $@������������������������       �                     @J       K                   ``@և���X�?             @������������������������       �                      @L       O                    �?���Q��?             @M       N                     Q@�q�q�?             @������������������������       �                      @������������������������       �                     �?P       Q                     Q@      �?              @������������������������       �                     �?������������������������       �                     �?S       X                   �Z@*T��Q�?�            �h@T       U                   �Y@؇���X�?             @������������������������       �                     @V       W                     J@�q�q�?             @������������������������       �                      @������������������������       �                     �?Y       l                   �j@D���"�?~            �g@Z       ]                    _@D�n�3�?#            �L@[       \                    �?$��m��?             :@������������������������       �                     1@������������������������       �                     "@^       g                   �h@��a�n`�?             ?@_       f                    @M@�eP*L��?             &@`       a                    �?      �?              @������������������������       �                     @b       c                   `h@���Q��?             @������������������������       �                     �?d       e                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @h       i                   @j@P���Q�?             4@������������������������       �                     *@j       k                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @m       �                   pn@�ʽ���?[            �`@n                           @P@�j��b�?&            �M@o       p                    �?@4և���?#             L@������������������������       �        	             *@q       v                   �_@�ʈD��?            �E@r       u                   pk@�nkK�?             7@s       t                   @k@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             2@w       z                   �`@R���Q�?             4@x       y                    �?      �?             @������������������������       �                      @������������������������       �                      @{       ~                   0k@      �?
             0@|       }                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@�       �                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   a@���+�?5            �R@�       �                    �?H(���o�?%            �J@�       �                    @O@      �?
             (@�       �                    �?�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?�4F����?            �D@������������������������       �        
             *@������������������������       �                     <@�       �                    �O@�����?             5@�       �                    �?�X�<ݺ?             2@������������������������       �                     �?������������������������       �                     1@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �e@l�;�	�?0            �R@�       �                    �?P�t��?/            @R@�       �                   Hs@8�A�0��?             6@�       �                    @Q@8�Z$���?             *@�       �                   �_@�8��8��?             (@�       �                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     "@������������������������       �                     �?�       �                   pu@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @�       �                    �?�\�u��?!            �I@������������������������       �                     0@������������������������       �                    �A@������������������������       �                      @�       �                   Xr@h8"J{�?[            �b@�       �                   l@�:�^���?R            �`@�       �                    �M@�IєX�?<            �Y@������������������������       �        "            �M@�       �                   �f@(L���?            �E@�       �                    �?"pc�
�?            �@@������������������������       �                     @������������������������       �                     ;@������������������������       �                     $@�       �                   �d@"pc�
�?            �@@�       �                    �M@      �?             8@�       �                   �o@�z�G��?             $@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �        	             ,@�       �                    �?�q�q�?             "@�       �                    �N@      �?             @������������������������       �                      @�       �                   �e@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   @u@      �?	             ,@�       �                    �?�<ݚ�?             "@�       �                    �J@�q�q�?             @������������������������       �                     �?�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h[�Bp       @a@     ��@     �]@      }@      V@     `z@      :@     @m@      :@      j@      0@      e@      *@      W@      &@     �V@      &@     �M@      @      &@       @      &@       @                      &@       @              @      H@       @      �?       @                      �?      @     �G@      @     �C@      @      5@       @      5@       @                      5@      �?                      2@       @       @      �?      @      �?       @               @      �?                      @      �?      �?      �?                      �?              @@       @      �?              �?       @              @     @S@              <@      @     �H@      �?               @     �H@              ,@       @     �A@              2@       @      1@       @                      1@      $@      D@      @      D@      @                      D@      @                      9@      O@     �g@      @      H@       @     �D@       @      B@              &@       @      9@       @       @              @       @       @      �?              �?       @      �?                       @              1@              @      @      @              @      @      @               @      @       @       @      �?       @                      �?      �?      �?              �?      �?             �L@     �a@      @      �?      @               @      �?       @                      �?     �I@     `a@      8@     �@@      1@      "@      1@                      "@      @      8@      @      @      @      @              @      @       @              �?      @      �?      @                      �?      @              �?      3@              *@      �?      @      �?                      @      ;@     �Z@      @     �J@      @      J@              *@      @     �C@      �?      6@      �?      @              @      �?                      2@      @      1@       @       @       @                       @      �?      .@      �?      @      �?                      @              (@       @      �?              �?       @              5@     �J@      3@      A@      @      @      @      @      @                      @      @              *@      <@      *@                      <@       @      3@      �?      1@      �?                      1@      �?       @      �?                       @      ?@      F@      =@      F@      *@      "@      &@       @      &@      �?       @      �?       @                      �?      "@                      �?       @      @              @       @              0@     �A@      0@                     �A@       @              3@     @`@      (@     �^@      @      X@             �M@      @     �B@      @      ;@      @                      ;@              $@      @      ;@      @      5@      @      @       @      �?              �?       @              �?      @      �?                      @              ,@      @      @      @      @       @              �?      @              @      �?                      @      @      @      @       @      @       @              �?      @      �?              �?      @              @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ	�tlhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvK)hwh(h+K ��h-��R�(KK)��h~�B�                            Xr@�Z{����?�           ��@                          �e@�����?�           Ѓ@                           �?�ftv���?j             d@������������������������       �        
             0@������������������������       �        `             b@       	                   @[@�Js
��?-           �}@                           �?�ՙ/�?             5@������������������������       �                     *@������������������������       �                      @
                           �J@=�AQ��?           @|@                           a@Ƶ�pD�?�             k@                           @B@����X�?]             d@������������������������       �                     "@                           �?|�i���?W             c@������������������������       �                     G@������������������������       �        =            �Z@                           �?4և����?$             L@������������������������       �                     @������������������������       �                     �I@                           �?X������?�            `m@������������������������       �                     A@������������������������       �        �             i@       (                     P@z�):���?8             Y@       #                    �J@�ݏ^���?2            �V@                            �?�!���?             A@                           �?���N8�?             5@������������������������       �                     �?                           �I@      �?             4@                           �?�n_Y�K�?	             *@������������������������       �                     @������������������������       �                      @������������������������       �                     @!       "                    �?��
ц��?             *@������������������������       �                     @������������������������       �                     @$       '                   {@      �?             L@%       &                    �?r�z-��?            �J@������������������������       �                    �A@������������������������       �        	             2@������������������������       �                     @������������������������       �                     $@�t�bh�h(h+K ��h-��R�(KK)KK��h[�B�        d@     ��@     �\@     @�@      0@      b@      0@                      b@     �X@     pw@      *@       @      *@                       @     @U@     �v@     �I@     �d@      G@     �\@              "@      G@     �Z@      G@                     �Z@      @     �I@      @                     �I@      A@      i@      A@                      i@      G@      K@      G@      F@      &@      7@      @      0@              �?      @      .@      @       @      @                       @              @      @      @      @                      @     �A@      5@     �A@      2@     �A@                      2@              @              $@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�ޡhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hK
hvKAhwh(h+K ��h-��R�(KKA��h~�B8                             �?�D����?�           ��@                           �?n\1�K��?�             w@                           �?Dc}h��?)             L@������������������������       �                     1@������������������������       �                    �C@                           �?��|��?�            �s@������������������������       �                     F@������������������������       �        �            �p@	       ,                    �?�W��0��?�            �v@
       +                   u@���h���?�            s@       (                   �`@�����?�            �r@                           �?v0���1�?x            `f@                          �Y@�����?g             c@                           @z�G�z�?             @                          �X@�q�q�?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           @�(�.Y��?c            `b@                           �?��k����?^             a@������������������������       �                    �E@������������������������       �        B            �W@                          �q@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?       '                    �L@X�<ݚ�?             ;@       &                   ``@���Q��?             9@       !                    @      �?             8@                            �?�E��ӭ�?             2@������������������������       �                     *@������������������������       �                     @"       %                   @_@�q�q�?             @#       $                   0l@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @)       *                    �?K�(i�?H            @]@������������������������       �                     3@������������������������       �        <            �X@������������������������       �                     "@-       <                    �?��.��?&            �N@.       9                   �q@d}h���?             E@/       6                    @K@�����H�?             B@0       5                    �J@�q�q�?             @1       2                   �`@z�G�z�?             @������������������������       �                      @3       4                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?7       8                    �?��S�ۿ?             >@������������������������       �                      @������������������������       �                     <@:       ;                   �b@r�q��?             @������������������������       �                     @������������������������       �                     �?=       @                    @I@�}�+r��?             3@>       ?                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        
             0@�t�bh�h(h+K ��h-��R�(KKAKK��h[�B       @d@     ��@     �N@     0s@      1@     �C@      1@                     �C@      F@     �p@      F@                     �p@     @Y@     �p@     �V@     �j@     �T@     �j@     �O@      ]@      H@      Z@      @      �?       @      �?      �?      �?      �?                      �?      �?               @              F@     �Y@     �E@     �W@     �E@                     �W@      �?      "@              "@      �?              .@      (@      .@      $@      .@      "@      *@      @      *@                      @       @      @       @      @       @                      @              �?              �?               @      3@     �X@      3@                     �X@      "@              $@     �I@      "@     �@@      @      @@       @      @      �?      @               @      �?       @      �?                       @      �?               @      <@       @                      <@      @      �?      @                      �?      �?      2@      �?       @      �?                       @              0@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJQY%hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hK	hvK;hwh(h+K ��h-��R�(KK;��h~�B�                              �?H�ig��?�           ��@                          Xr@���ɕ��?�            �x@                           �N@�.nq�?�            u@                           �?țu���?�            @p@������������������������       �                     ;@������������������������       �        �             m@                           [@��مD�?0            @S@������������������������       �                     @	       
                    �?��G���?.            �R@������������������������       �                     ,@������������������������       �        &             N@                          �t@:2vz�M�?%            �N@                            P@ҳ�wY;�?             A@                          �r@>���Rp�?             =@                           �?      �?              @������������������������       �                     @������������������������       �                     @                           �?�����?	             5@������������������������       �                     3@������������������������       �                      @������������������������       �                     @                           �?PN��T'�?             ;@                          �`@      �?             @������������������������       �                     �?������������������������       �                     @                           �?�nkK�?             7@                           b@      �?             0@������������������������       �                     &@                           �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @!       $                    �?�q�q�?�             u@"       #                    �?����b�?�             q@������������������������       �        7            @V@������������������������       �        ~             g@%       :                    �?���-T��?'             O@&       +                    `@��P���?            �D@'       (                    @      �?             0@������������������������       �                     *@)       *                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?,       9                     Q@ �o_��?             9@-       8                    �L@��<b���?             7@.       3                   k@X�Cc�?             ,@/       0                   �h@      �?              @������������������������       �                     @1       2                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?4       5                    �?�q�q�?             @������������������������       �                      @6       7                   �`@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     "@������������������������       �                      @������������������������       �                     5@�t�bh�h(h+K ��h-��R�(KK;KK��h[�B�        e@     ��@     �Q@     �t@      F@     Pr@      ;@      m@      ;@                      m@      1@      N@      @              ,@      N@      ,@                      N@      :@     �A@      6@      (@      6@      @      @      @      @                      @      3@       @      3@                       @              @      @      7@      @      �?              �?      @              �?      6@      �?      .@              &@      �?      @      �?                      @              @     �X@     �m@     @V@      g@     @V@                      g@      "@     �J@      "@      @@       @      ,@              *@       @      �?       @                      �?      @      2@      @      2@      @      "@      �?      @              @      �?       @               @      �?              @       @       @               @       @       @                       @              "@       @                      5@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��fbhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hK
hvKhwh(h+K ��h-��R�(KK��h~�B�                            Xr@�6�L���?�           ��@                           �?�@�����?�           �@������������������������       �        J            �\@������������������������       �        N           X�@                           @F@�d�~V��?;            @X@������������������������       �        	             .@                           �?z�^��?2            �T@                           @O@��C���?            �G@	                          �t@�Q����?             D@
                          �_@��H�}�?             9@������������������������       �                      @                           �?8����?             7@                          @s@b�2�tk�?
             2@                           �N@������?             .@                           �?d}h���?             ,@������������������������       �                     &@������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                           �?z�G�z�?             .@������������������������       �                     @������������������������       �        	             (@������������������������       �                     @                           �?��R[s�?            �A@������������������������       �                     :@������������������������       �                     "@�t�bh�h(h+K ��h-��R�(KKKK��h[�B�       �c@     ��@     �\@     X�@     �\@                     X�@     �F@      J@              .@     �F@     �B@      3@      <@      3@      5@      0@      "@               @      0@      @      &@      @      &@      @      &@      @      &@                      @              �?              @      @              @      (@      @                      (@              @      :@      "@      :@                      "@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ$�phG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvKhwh(h+K ��h-��R�(KK��h~�B                             �?�`��ie�?�           ��@                          l@L)Þ\��?�            �x@                           �?L���
B�?~            �i@������������������������       �                     0@������������������������       �        q            �g@                           �?�YT�� �?l            `g@������������������������       �                    �C@������������������������       �        U            �b@	                          �p@Dn����?�            @u@
                           �?"pc�
�?�            �p@������������������������       �        $             H@������������������������       �        }             k@                          �_@��}�+r�?3             S@                           @B@�<ݚ�?             ;@������������������������       �                      @                           �?�J�4�?             9@������������������������       �                     5@������������������������       �                     @                           �G@Tt�ó��?"            �H@������������������������       �                     &@                           �?D�n�3�?             C@������������������������       �                     6@������������������������       �                     0@�t�bh�h(h+K ��h-��R�(KKKK��h[�Bp       @b@     `�@     �K@     0u@      0@     �g@      0@                     �g@     �C@     �b@     �C@                     �b@     �V@      o@      H@      k@      H@                      k@     �E@     �@@      5@      @               @      5@      @      5@                      @      6@      ;@              &@      6@      0@      6@                      0@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJW:+LhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvKhwh(h+K ��h-��R�(KK��h~�C�                           �?N8���?�           ��@������������������������       �        j            @e@������������������������       �        l           ��@�t�bh�h(h+K ��h-��R�(KKKK��h[�C0     @e@     ��@     @e@                     ��@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJF<KdhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvK?hwh(h+K ��h-��R�(KK?��h~�B�         .                    �?$r�%oR�?�           ��@       +                   �b@������?�            �v@                           �?��8���?�            �q@                           �?l��w��?�            �i@                          Pm@���c���?$             J@������������������������       �                     6@                          �_@�������?             >@                          p@$�q-�?             *@	       
                   `o@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@                          o@ҳ�wY;�?             1@������������������������       �                      @                          Xp@������?
             .@������������������������       �                     @                          �`@���Q��?             $@                          �s@      �?             @������������������������       �                     @������������������������       �                     �?                          �r@r�q��?             @������������������������       �                     @                          b@      �?              @������������������������       �                     �?������������������������       �                     �?                           �?��T��g�?e            @c@������������������������       �                     9@������������������������       �        V             `@       (                   �t@ףp=
�?.             T@       '                    �?@-�_ .�?,            �R@       "                   `Z@l�b�G��?"            �L@        !                    �?���!pc�?             &@������������������������       �                     @������������������������       �                      @#       &                   �\@��<b�ƥ?             G@$       %                    \@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                    �B@������������������������       �        
             1@)       *                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @,       -                    �?�d�����?4             S@������������������������       �                     4@������������������������       �        '             L@/       >                   �u@4�S�#W�?�            @w@0       ;                    f@�� -!��?�            �v@1       6                    �?     p�?%             P@2       5                    @F@ "��u�?             I@3       4                    �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     F@7       :                    �?؇���X�?             ,@8       9                    @�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     @<       =                    �?������?�            �r@������������������������       �        9            @U@������������������������       �        �            @k@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK?KK��h[�B�       `c@     �@      N@     �r@      D@     �n@      @@     �e@      @     �F@              6@      @      7@      �?      (@      �?      @              @      �?                      "@      @      &@       @              @      &@              @      @      @      @      �?      @                      �?      �?      @              @      �?      �?              �?      �?              9@      `@      9@                      `@       @      R@      @     �Q@      @     �J@      @       @      @                       @      �?     �F@      �?       @               @      �?                     �B@              1@      @       @               @      @              4@      L@      4@                      L@     �W@     Pq@     �V@     Pq@      @     �M@      @     �G@      @      @      @                      @              F@       @      (@       @      @              @       @                      @     @U@     @k@     @U@                     @k@      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJؽ�hG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hK	hvKGhwh(h+K ��h-��R�(KKG��h~�B�         (                    @K@D�w@B��?�           ��@                          �h@�z�G��?�            �w@                           �D@���c���?A             Z@                           �?">�֕�?            �A@                           �?�5��?             ;@                          �e@�d�����?             3@       
                    �C@8�Z$���?	             *@       	                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     "@                           �?      �?             @������������������������       �                     @������������������������       �                     @                          Pb@      �?              @������������������������       �                     �?                           @C@؇���X�?             @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @                          �c@�nkK�?+            @Q@                           �?Pa�	�?(            �P@������������������������       �                      @������������������������       �        &             P@                           �?�q�q�?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?        #                    �?�#��ؒ�?�            @q@!       "                    �?�^����?�            @n@������������������������       �        +            �T@������������������������       �        g            �c@$       '                    b@      �?             A@%       &                    �?��}*_��?             ;@������������������������       �                     1@������������������������       �                     $@������������������������       �                     @)       @                    �?�k�#��?�             v@*       -                    �?�4���L�?�             p@+       ,                    �?�՘���?x            �g@������������������������       �                     F@������������������������       �        ]            @b@.       ;                   �l@ДX��?/             Q@/       0                    �?�r����?            �F@������������������������       �                     *@1       :                   @l@     ��?             @@2       5                   �Y@�r����?             >@3       4                    @N@      �?             @������������������������       �                     �?������������������������       �                     @6       7                    c@ ��WV�?             :@������������������������       �                     1@8       9                    �?�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                      @<       =                   Hr@�nkK�?             7@������������������������       �                     0@>       ?                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @A       D                   Pr@�8��8N�?>             X@B       C                    �?��+��<�?7            �U@������������������������       �                     @������������������������       �        4            �T@E       F                    �?���Q��?             $@������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KKGKK��h[�Bp       �e@     ��@     �\@     �p@      ,@     �V@      &@      8@      &@      0@      @      ,@       @      &@       @       @       @                       @              "@      @      @              @      @              @       @              �?      @      �?       @      �?       @                      �?      @                       @      @     �P@       @      P@       @                      P@      �?       @      �?      �?              �?      �?                      �?      Y@      f@     �T@     �c@     �T@                     �c@      1@      1@      1@      $@      1@                      $@              @      M@     �r@     �I@     �i@      F@     @b@      F@                     @b@      @     �N@      @     �C@              *@      @      :@      @      :@      @      �?              �?      @              �?      9@              1@      �?       @      �?                       @       @              �?      6@              0@      �?      @      �?                      @      @     @V@      @     �T@      @                     �T@      @      @      @                      @�t�bub��      hhubh)��}�(hhhhhNhKhKhG        hh$hNhJX��vhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvKhwh(h+K ��h-��R�(KK��h~�C�                           �?�'�Ռ��?�           ��@������������������������       �        h             e@������������������������       �        i           ��@�t�bh�h(h+K ��h-��R�(KKKK��h[�C0      e@     ��@      e@                     ��@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���EhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvKhwh(h+K ��h-��R�(KK��h~�Bh                             s@�6�L���?�           ��@                           �?����?�           ��@������������������������       �        T            �_@������������������������       �        Q           ��@                           �?      �?+            �P@                           �?��S���?'             N@������������������������       �                     @@������������������������       �                     <@	       
                   `@r�q��?             @������������������������       �                     �?������������������������       �                     @�t�bh�h(h+K ��h-��R�(KKKK��h[�C�     �c@     ��@     �_@     ��@     �_@                     ��@     �@@     �@@      @@      <@      @@                      <@      �?      @      �?                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ:9)bhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvK9hwh(h+K ��h-��R�(KK9��h~�Bx         8                   �h@>��g/�?�           ��@       5                    @K@��a1��?�           ��@                            �?Pu�����?�             x@                          `a@r�,����?q            @f@                          0m@R�c���?O             `@                          �`@�5U��K�?2            �T@                           �I@ĴF���?1            �T@                          �[@�]0��<�?$            �N@	                           �G@���}<S�?             7@
                          @M@���N8�?             5@                           �?      �?              @                           �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     *@                          `T@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     C@                           `@���N8�?             5@������������������������       �        	             (@                          �V@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     �?                           �?\X��t�?             G@������������������������       �                     4@������������������������       �                     :@                           �?@9G��?"            �H@������������������������       �                      @������������������������       �                     �G@!       2                    @I@���3�E�?{             j@"       /                    �?�tk~X$�?W             b@#       ,                   �`@�v:���?.             Q@$       +                    �?      �?#             H@%       (                    @E@
;&����?"             G@&       '                    �?l��
I��?             ;@������������������������       �                      @������������������������       �                     3@)       *                    �?�d�����?             3@������������������������       �                     ,@������������������������       �                     @������������������������       �                      @-       .                   @r@P���Q�?             4@������������������������       �        
             3@������������������������       �                     �?0       1                    �?p9W��S�?)             S@������������������������       �                     6@������������������������       �                     K@3       4                    �?     ��?$             P@������������������������       �        	             *@������������������������       �                    �I@6       7                    �?N���X�?�            �u@������������������������       �        &             J@������������������������       �        �            `r@������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK9KK��h[�B�        b@     p�@     �a@     p�@     �V@     �r@      >@     �b@      <@     @Y@       @     �R@      @     �R@       @     �M@       @      5@      �?      4@      �?      @      �?      @      �?                      @              @              *@      �?      �?              �?      �?                      C@      @      0@              (@      @      @              @      @              �?              4@      :@      4@                      :@       @     �G@       @                     �G@      N@     �b@     �G@     @X@      9@     �E@      8@      8@      6@      8@       @      3@       @                      3@      ,@      @      ,@                      @       @              �?      3@              3@      �?              6@      K@      6@                      K@      *@     �I@      *@                     �I@      J@     `r@      J@                     `r@       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�BHzhG        hNhG        hAKhBKhCh(h+K ��h-��R�(KK��h[�C              �?�t�bhOh`hcC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hc�C       �t�bK��R�}�(hKhvKhwh(h+K ��h-��R�(KK��h~�Bh                            �e@��Mw��?�           ��@                           �?�Z<p���?�           0�@������������������������       �        W             a@������������������������       �        b           �@       
                   0r@r�q��?             8@       	                   `f@     ��?
             0@                          �\@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@������������������������       �                      @�t�bh�h(h+K ��h-��R�(KKKK��h[�C�     �b@     P�@      a@     �@      a@                     �@      &@      *@      @      *@      @      �?              �?      @                      (@       @        �t�bubhhubehhub.